!!!! CIURCUIT !!!!
V1VAR n1 0 PWL(0 0 1e-9 0)
R1 n2 n1 {parR1}
C1 n2 0 {parC1}
.param parR1=100
.param parC1=500e-6
.ic V(n1)=0
**********MODELS**********
*****MODEL1*****
